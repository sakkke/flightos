module main

const default_config_map = {
	'console_keymap': ['us']
	'disk':           ['/dev/sda']
}
