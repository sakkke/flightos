module main

const default_config_map = {
	'console_keymap':    ['us']
	'disk':              ['/dev/sda']
	'installation_mode': ['Custom']
	'locale':            ['en_US.UTF-8 UTF-8']
	'packages':          []
	'timezone':          ['UTC']
}
